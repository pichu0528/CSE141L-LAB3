import definitions::*;

// This a simple memory module which simulates the cache for the core, with handshake features. 
// Handshake method description: the core sends a request for read or write (valid signal). 
// Memory responses in time (yumi signal).
// Memory sends the valid signal afterwards and the required data if any. 
// Finally memory waits for the core until it receives the yumi signal from the core. 
// Input and output structures are defined in definitions.v file
// IDLE means the memory is waiting for a request. TRANS means the memory 
// is during a data transaction and it is waiting for the core to response yumi.

module data_mem #(
        parameter addr_width_p = 12
    )
    (
        input  clk,
        input  n_reset,
        input  [$bits(mem_in_s)-1:0]  port_flat_i,
        input  [31:0] addr,     // we accept a 32-bit address
        output [$bits(mem_out_s)-1:0] port_flat_o
    ); 

    // Flatten and Unflatten structs
    mem_in_s port_i;
    mem_out_s port_o;
    assign port_i = port_flat_i;
    assign port_flat_o = port_o;

    logic [7:0] mem [(2**addr_width_p)-1];

    //Registers
    logic wen_r;
    logic [31:0] read_data_r;

    enum logic{
        IDLE  = 1'b0,
        TRANS = 1'b1
    } state_r;

    logic port_i_wen_override;

    // don't write if the address is out of bounds
    assign port_i_wen_override = port_i.wen & ~|(addr >> addr_width_p);

    always_ff @ (negedge clk)
        begin
        if (~port_i.byte_not_word & (| addr[1:0]) & port_i_wen_override)
            begin
            $display("ERROR: unaligned word write of data %x to address %x\n",port_i.write_data, addr);
        end
    end
  

    always_ff @ (posedge clk)
    begin
        port_o.valid     <= 1'b0;
        port_o.read_data <= 32'bx;
        read_data_r      <= 32'bx;
        if (!n_reset)
            begin
            state_r      <= IDLE;
            end
        else
            begin
            unique case (state_r)
                IDLE:
                    begin
                    if (port_i.valid) 
                        begin        
                        state_r      <= TRANS;
                        port_o.valid <= 1'b1;
                        
                        // mbt: don't write if address out of bounds
                        wen_r   <= port_i_wen_override;
                        if (port_i_wen_override)
                            begin
                            if (port_i.byte_not_word)
                                begin
                                mem [addr] <= port_i.write_data[7:0];
                                end
                            else
                                begin
                                {mem[addr+3],mem[addr+2],mem[addr+1],mem[addr]}<=port_i.write_data;
                            end
                            end
                        else
                            begin   
                            if (port_i.byte_not_word)
                                begin
                                port_o.read_data <= {{24{1'b0}}, {mem[addr]}};
                                read_data_r      <= {{24{1'b0}}, {mem[addr]}};
                                end
                            else
                                begin
                                port_o.read_data <= {mem[addr+3], mem[addr+2], mem[addr+1], mem[addr]};
                                read_data_r      <= {mem[addr+3], mem[addr+2], mem[addr+1], mem[addr]};
                            end
                        end
                        end // if
                    else
                        begin
                        state_r <= IDLE;
                    end
                end
                
                TRANS:
                    begin
                    if (port_i.yumi)
                        begin
                        state_r        <= IDLE;
                        end
                    else
                        begin
                        port_o.valid <= 1'b1;
                        state_r      <= TRANS;
                        wen_r        <= wen_r;
                        read_data_r  <= read_data_r;
                        if (!wen_r)
                            begin
                            port_o.read_data <= read_data_r;
                        end
                    end
                end
                    
                default:
                    state_r <= IDLE;

            endcase
        end
    end

    // Since there is no delay for this memory, as soon as it gets the valid signal from 
    // the core memory responses yumi which means I recieved the signal, and data in store mode.
    always_comb
        begin
        port_o.yumi = port_i.valid;
    end

endmodule
